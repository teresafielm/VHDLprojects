library IEEE; --Librerías
use IEEE.STD_LOGIC_1164.ALL; --Liberías
ENTITY Deco is --Definimos entidad
PORT ( Q,W,E,R,T,Y,U,I: in STD_LOGIC; X,IC,S,A,O,N,C,J,RE,M,D : out STD_LOGIC); 
--Decodificador de 8 entradas y 11 salidas
END Deco; --Se termina entidad
ARCHITECTURE Behavioral OF Deco IS --Iniciamos arquitectura
BEGIN
X<= NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND NOT Y AND 
NOT U AND NOT I; --XOR--
IC<=NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND NOT Y AND 
NOT U AND I;-- INVERTIR--
S<= NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND NOT Y AND U 
AND NOT I;--SUMA--
A<= NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND NOT Y AND U 
AND I;--AND--
O<= NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND Y AND NOT U 
AND NOT I;--OR--
N<= NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND Y AND NOT U 
AND I ;--NO OPERACIÓN--
C<= NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND Y AND U AND 
NOT I;--CARGA--
J<= NOT Q AND NOT W AND NOT E AND NOT R AND NOT T AND Y AND U AND 
I;--JUMP--
RE<=NOT Q AND NOT W AND NOT E AND NOT R AND T AND NOT Y AND NOT U 
AND NOT I ;--RESTA--
M<= NOT Q AND NOT W AND NOT E AND NOT R AND T AND NOT Y AND NOT U 
AND I ;--MULTIIPLICACIÓN--
D<= NOT Q AND NOT W AND NOT E AND NOT R AND T AND NOT Y AND U AND 
NOT I;--DIVISIÓN--
END Behavioral; --Final de arquitectura